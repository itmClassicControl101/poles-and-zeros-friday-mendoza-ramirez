;LC circuit for space-states:
;Vin 1 0 pulse (0.5, 5V, 0s, 1ns, 1ns, 1ms, 2ms)
Vin 1 0 AC 5
R1 1 2 10k
R2 2 3 10k
R3 2 0 10k
L1 3 0 4.25mF
;.tran 100us 4ms
.ac dec 10 10Hz 100000k
.probe
.end